library IEEE;
use IEEE.std_logic_1164.all;

entity completeMDR is
port(
something : IN std_logic
);

architecture behavior of muxMDR is
BEGIN

END architecture;